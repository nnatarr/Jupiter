��- - - - - - - - - - - - - - - - - - - - -   C e l l   m y C e l l   - - - - - - - - - - - - - - - - - - - - - -  
 e n t i t y   m y C e l l   i s   p o r t ( x 0 ,   x 1 ,   x 2 ,   x 3 :   i n   B I T ;   y :   o u t   B I T ) ;  
     e n d   m y C e l l ;  
  
 a r c h i t e c t u r e   m y C e l l _ B O D Y   o f   m y C e l l                   i s  
     c o m p o n e n t   2 b a n d 2 _ o r 2   p o r t ( X 1 ,   X 2 ,   X 3 ,   X 4 :   i n   B I T ;   Z :   o u t   B I T ) ;  
         e n d   c o m p o n e n t ;  
  
     s i g n a l   i n v _ 0 ,   i n v _ 1 ,   i n v _ 2 ,   n e t _ 0 ,   n e t _ 1 :   B I T ;  
  
 b e g i n  
     E L M 2 :   2 b a n d 2 _ o r 2   p o r t   m a p ( i n v _ 1 ,   n e t _ 0 ,   x 1 ,   n e t _ 1 ,   y ) ;  
     E L M 1 :   2 b a n d 2 _ o r 2   p o r t   m a p ( i n v _ 0 ,   0 ,   0 ,   x 2 ,   n e t _ 1 ) ;  
     E L M 0 :   2 b a n d 2 _ o r 2   p o r t   m a p ( i n v _ 2 ,   0 ,   0 ,   i n v _ 0 ,   n e t _ 0 ) ;  
     P S E U D O _ I N V E R T 2 :   i n v e r t e r   p o r t   m a p ( x 3 ,   i n v _ 2 ) ;  
     P S E U D O _ I N V E R T 1 :   i n v e r t e r   p o r t   m a p ( x 1 ,   i n v _ 1 ) ;  
     P S E U D O _ I N V E R T 0 :   i n v e r t e r   p o r t   m a p ( x 0 ,   i n v _ 0 ) ;  
 e n d   m y C e l l _ B O D Y ; 